module mux4_1_tb();

  reg [1:0]sel;
  reg [3:0]a;
  wire y ;

  integer i,j;
// Instantiate the Design 
  mux4_1 DUT(.a(a), .sel(sel), .y(y));

  task initialize;
  begin 
		a=0;
    sel=0;
  end
  endtask

  task select(input [1:0]s);
  begin
    sel=s;
  end
  endtask
 
  task inps(input[3:0] data);
  begin
    a=data;
  end
  endtask

initial 
begin
  initialize;
  #10;
  for(i=0;i<4;i=i+1)
  begin
    select(i);
    for(j=0;j<16;j=j+1)
    begin
      inps(j);
      #10;
    end
  end
end
// Use $monitor task in a parallel initial block  to display inputs and outputs.

initial 
  $monitor("a[3:0]=%b--select=%b--y=%d\n",a,sel,y);

// Use $finish task to finish the simulation in a parallel initial block with appropriate delay.
initial 

#800 $finish;

endmodule